LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY P7194 IS
PORT(V : IN STD_LOGIC_VECTOR(3 downto 0);
     CLK, CLR, S0, S1, SR, SL : IN STD_LOGIC;
     Q: OUT STD_LOGIC_VECTOR(3 downto 0));
END P7194;

ARCHITECTURE BEHAVIORAL OF P7194 IS
SIGNAL G,QA: STD_LOGIC_VECTOR(3 downto 0);
BEGIN
G <= QA;
PROCESS(CLK,CLR)
BEGIN
IF (CLR = '0') THEN
QA <= "0000";
ELSIF (rising_edge(CLK)) THEN
IF (S0 = '1' and S1 = '1') THEN
QA <= V;
ELSIF (S0 = '0' and S1 = '1') THEN
QA <= SR & G(3 downto 1);
ELSIF (S0 = '1' and S1 = '0') THEN QA <= G(2 downto 0) & SL;
ELSIF (S0 = '0' and S1 = '0') THEN
QA <= QA;
END IF;
END IF;
Q <= QA;
END PROCESS;
END BEHAVIORAL;
