LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY EJ1 IS
PORT(VE: IN STD_LOGIC_VECTOR(7 downto 0);
     VS: OUT STD_LOGIC_VECTOR(7 downto 0);
     CLKB, CLRB, S0B, S1B: in STD_LOGIC);
end EJ1;

ARCHITECTURE BEHAVIORAL OF EJ1 IS
COMPONENT P7194
PORT (V : IN STD_LOGIC_VECTOR(3 downto 0);
     CLK, CLR, S0, S1, SR, SL : IN STD_LOGIC;
     Q: OUT STD_LOGIC_VECTOR(3 downto 0));
END COMPONENT;

SIGNAL ACT: STD_LOGIC_VECTOR(7 downto 0):= "00000000";
BEGIN
VS <= ACT;
P0: P7194 PORT MAP(VE(7 downto 4), CLKB, CLRB, S0B, S1B, ACT(3), ACT(0), ACT(7 downto 4));
P1: P7194 PORT MAP(VE(3 downto 0), CLKB, CLRB, S0B, S1B, ACT(7), ACT(4), ACT(3 downto 0));
END BEHAVIORAL;
