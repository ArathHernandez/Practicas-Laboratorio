LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY P74F169 is
port ( UD, CLK1, CEP, CET, PE : IN STD_LOGIC;
D : IN STD_LOGIC_VECTOR( 3 downto 0);
Q : OUT STD_LOGIC_VECTOR (3 downto 0);
TC: OUT STD_LOGIC);
END P74F169;

ARCHITECTURE BEHAVIORAL OF P74F169 IS
SIGNAL t: STD_LOGIC_VECTOR(3 downto 0):="0000";
SIGNAL r: STD_LOGIC := '1';
BEGIN
TC <= r;
PROCESS(CLK1, r, PE)
BEGIN
IF (CET = '0' and CEP = '0') THEN
IF(rising_edge(CLK1))THEN
IF(UD = '1')THEN
t <= t+1;
IF (t = "1001") THEN
t <= "0000";
r <= '0';
ELSE
r <= '1';
END IF;
ELSE
t <= t-1;
IF (t = "0000") THEN
t <= "1001";
r <= '0';
ELSE
r <= '1';
END IF;
END IF;
END IF;
IF (PE = '0') THEN
t <= D;
END IF;
END IF;
END PROCESS;
Q <= t;
END BEHAVIORAL;
